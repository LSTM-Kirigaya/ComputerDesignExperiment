`include "./DataPath/alu_ctrl.v"
`include "./DataPath/alu.v"
`include "./DataPath/dm.v"
`include "./DataPath/Ext.v"
`include "./DataPath/im.v"
`include "./DataPath/mux.v"
`include "./DataPath/npc.v"
`include "./DataPath/pc.v"
`include "./DataPath/pc_add.v"
`include "./DataPath/regfile.v"
`include "./DataPath/branch_add.v"
`include "./DataPath/IF_ID.v"
`include "./DataPath/ID_EX.v"
`include "./DataPath/EX_MEM.v"
`include "./DataPath/MEM_WB.v"

module data_path(
    LS_bit,
    RegDst, 
    Branch, 
    MemtoReg, 
    ALUOp, 
    MemWrite, 
    ALUSrc, 
    RegWrite, 
    Jump, 
    Ext_op, 
    PctoReg,

    clock, 
    reset,

    IF_ID_out
    
    );

    input   [ 1: 0] LS_bit;
    input           RegDst;
    input   [ 1: 0] Branch;
    input           MemtoReg;
    input   [ 3: 0] ALUOp;
    input           MemWrite;
    input           ALUSrc;
    input           RegWrite;
    input           Jump;
    input           Ext_op;
    input           PctoReg;

    input           clock;
    input           reset;

    output  [63: 0] IF_ID_out;

    // variable
    wire    [31: 0] PC;             // value of pc
    wire    [31: 0] NPC;            // next status of pc 
    wire    [31: 0] ext_out;        // extention of 16-bit   
    wire    [31: 0] instruction;    // instruction gotten by im
    wire            zero;           // zero generated by ALU
    wire    [31: 0] pc_add_out;     // pc + 4

    wire    [31: 0] regfile_out1;   // out1 of regfile
    wire    [31: 0] regfile_out2;   // out2 of regfile

    wire    [ 4: 0] mux1_out;       // IF ID
    wire    [31: 0] mux2_out;       // ID EX
    wire    [31: 0] mux3_out;       // MEM WB
    wire    [31: 0] mux4_out;
    wire    [ 4: 0] mux5_out;
    wire    [31: 0] mux6_out;

    wire    [ 3: 0] alu_ctrl_out;   // out of alu controller
    wire    [31: 0] alu_out;        // out of alu
    wire    [31: 0] dm_out;         // out of dm
    wire    [31: 0] branch_add_out; // out of branch add

    // pipeline register
    wire    [63 : 0] IF_ID_out;
    wire    [137: 0] ID_EX_out;
    wire    [169: 0] EX_MEM_out;
    wire    [103: 0] MEM_WB_out;

    // pc module
    pc program_counter(
        .NPC(NPC),
        .clock(clock),
        .reset(reset),
        .PC(PC)
    );

    pc_add pc_adder(
        .PC(PC),
        .pc_add_out(pc_add_out)
    );

    npc next_program_counter(
        .Jump(Jump),
        .branch(Branch),
        .zero(zero),
        .EX_MEM_branch_add_out(EX_MEM_out[40:9]),
        .EX_MEM_pc_add_out(EX_MEM_out[73:42]),
        .EX_MEM_instr26(EX_MEM_out[99:74]),
        .NPC(NPC)
    );

    // IF module, from pc value to the cycle's instructions
    im_4k instruction_memory(
        .pc(PC),
        .out_instr(instruction)
    );

    // IF/ID 
    IF_ID IF_ID_pipeline_register(
        .clock(clock),
        .pc_add_out(pc_add_out),
        .im_out(instruction),
        .IF_ID_out(IF_ID_out)
    );

    // ID module
    regfile register_files(
        .rs(IF_ID_out[57:53]),
        .rt(IF_ID_out[52:48]),
        .rd(mux5_out),
        .data(mux4_out),
        .RegWrite(MEM_WB_out[0]),
        .clock(clock),
        .reset(reset),
        .regfile_out1(regfile_out1),
        .regfile_out2(regfile_out2)
    );

    // ID/EX
    ID_EX ID_EX_pipeline_register(
        .clock(clock),
        .reset(reset),

        .LS_bit(LS_bit),
        .RegDst(RegDst),
        .Branch(Branch),
        .MemtoReg(MemtoReg),
        .ALUOp(ALUOp),
        .MemWrite(MemWrite),
        .Jump(Jump),
        .Ext_op(Ext_op),
        .PctoReg(PctoReg),
        
        .IF_ID_pc_add_out(IF_ID_out[31:0]),
        .regfile_out1(regfile_out1),
        .regfile_out2(regfile_out2),
        .instr26(IF_ID_out[57:32]),

        .ID_EX_out(ID_EX_out)
    );

    // EX module
    mux1 u_mux1(
        .rt(ID_EX_out[132:128]),
        .rd(ID_EX_out[127:123]),
        .RegDst(ID_EX_out[2]),
        .DstReg(mux1_out)
    );

    Ext extension_unit(
        .input_num(ID_EX_out[127:112]),
        .Ext_op(ID_EX_out[14]),
        .output_num(ext_out) 
    );

    alu_ctrl ALU_controller(
        .funct(ext_out[5:0]),           // last 5 bit of instruction, which repersents funct code
        .ALUOp(ID_EX_out[9:6]),         // ALUOp
        .alu_ctrl_out(alu_ctrl_out)
    );

    mux2 u_mux2(
        .out2(ID_EX_out[111:80]),        // regfile_out2
        .Ext(ext_out),
        .ALUSrc(ID_EX_out[11]),          // ALUSrc
        .DstData(mux2_out)
    );

    alu ALU(
        .op_num1(ID_EX_out[79:48]),     // regfile_out1
        .op_num2(mux2_out),
        .shamt(ext_out[10:6]),  
        .alu_ctrl_out(alu_ctrl_out),
        .zero(zero),
        .alu_out(alu_out)
    );

    branch_add branch_move_adder(
        .ID_EX_pc_add_out(ID_EX_out[47:16]),
        .Ext_out(ext_out),
        .branch_add_out(branch_add_out)
    );

    mux6 u_mux6(
        .ID_EX_pc_add_out(ID_EX_out[47:16]),
        .ID_EX_regfile_out2(ID_EX_out[111:80]),
        .funct(ID_EX_out[117:112]),
        .mux6_out(mux6_out)
    );  


    // EX/MEM
    EX_MEM EX_MEM_pipeline_register(
        .clock(clock),
        .reset(reset),

        .LS_bit(LS_bit),
        .Branch(ID_EX_out[4:3]),
        .MemtoReg(ID_EX_out[5]),
        .MemWrite(ID_EX_out[10]),
        .RegWrite(ID_EX_out[12]),
        .Jump(ID_EX_out[13]),
        .Ext_op(ID_EX_out[14]),
        .PctoReg(ID_EX_out[15]),

        .branch_add_out(branch_add_out),
        .zero(zero),
        .ID_EX_pc_add_out(mux6_out),
        .ID_EX_instr26(ID_EX_out[137:112]),
        .alu_out(alu_out),
        .ID_EX_regfile_out2(ID_EX_out[111:80]),
        .mux1_out(mux1_out),

        .EX_MEM_out(EX_MEM_out)
    );

    
    // MEM module
    dm_4k data_memory(
        .clock(clock),
        .EX_MEM_alu_out(EX_MEM_out[132:101]),
        .EX_MEM_register_out2(EX_MEM_out[164:133]),
        .LS_bit(EX_MEM_out[1:0]),
        .MemWrite(EX_MEM_out[2]),
        .Ext_op(EX_MEM_out[8]),
        .dm_out(dm_out)
    );

    // MEM/WB
    MEM_WB MEM_WB_pipeline_register(
        .clock(clock),
        .reset(reset),

        .RegWrite(EX_MEM_out[6]),
        .MemtoReg(EX_MEM_out[4]),
        .PctoReg(EX_MEM_out[9]),

        .EX_MEM_pc_add_out(EX_MEM_out[74:43]),
        .dm_out(dm_out),
        .EX_MEM_alu_out(EX_MEM_out[132:101]),
        .EX_MEM_mux1_out(EX_MEM_out[169:165]),

        .MEM_WB_out(MEM_WB_out)
    );

    // WB module
    mux3 u_mux3(
        .dm_out(MEM_WB_out[66:35]),
        .alu_out(MEM_WB_out[98:67]),
        .MemtoReg(MEM_WB_out[1]),
        .mux3_out(mux3_out)
    );


    mux4 u_mux4(
        .mux3_out(mux3_out),
        .MEM_WB_pc_add_out(MEM_WB_out[34:3]),
        .PctoReg(MEM_WB_out[2]),
        .mux4_out(mux4_out)
    );

    mux5 u_mux5(
        .MEM_WB_mux1_out(),
        .PctoReg(),
        .mux5_out(mux5_out)
    );

endmodule
