module HDU1 (
    input    [ 4: 0] rs,
    input    [ 4: 0] rt,
    input    [ 4: 0] mux1_out

);

endmodule // HDU1

module HDU2 (
    
);

endmodule //HDU2