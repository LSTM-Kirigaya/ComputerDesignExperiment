module v3();
    initial begin
        $display("I am v3");
    end
endmodule //v3