module datapath (
    
);

endmodule //datapath