module EPC (
    
);

endmodule //EPC