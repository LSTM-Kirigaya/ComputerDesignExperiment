`include "./DataPath/alu_ctrl.v"
`include "./DataPath/alu.v"
`include "./DataPath/dm.v"
`include "./DataPath/Ext.v"
`include "./DataPath/im.v"
`include "./DataPath/mux.v"
`include "./DataPath/npc.v"
`include "./DataPath/pc.v"
`include "./DataPath/pc_add.v"
`include "./DataPath/regfile.v"
`include "./DataPath/branch_add.v"
`include "./DataPath/IF_ID.v"
`include "./DataPath/ID_EX.v"
`include "./DataPath/EX_MEM.v"
`include "./DataPath/MEM_WB.v"

module data_path(
    LS_bit,
    RegDst, 
    Branch, 
    MemtoReg, 
    ALUOp, 
    MemWrite, 
    ALUSrc, 
    RegWrite, 
    Jump, 
    Ext_op, 
    PctoReg,

    clock, 
    reset,

    IF_ID_im_out
    
    );

    input   [ 1: 0] LS_bit;
    input           RegDst;
    input   [ 1: 0] Branch;
    input           MemtoReg;
    input   [ 3: 0] ALUOp;
    input           MemWrite;
    input           ALUSrc;
    input           RegWrite;
    input           Jump;
    input           Ext_op;
    input           PctoReg;

    input           clock;
    input           reset;

    output  [31: 0] IF_ID_im_out;


    // variable
    wire    [31: 0] PC;             // value of pc
    wire    [31: 0] NPC;            // next status of pc 
    wire    [31: 0] ext_out;        // extention of 16-bit   
    wire    [31: 0] instruction;    // instruction gotten by im
    wire            zero;           // zero generated by ALU
    wire    [31: 0] pc_add_out;     // pc + 4

    wire    [31: 0] regfile_out1;   // out1 of regfile
    wire    [31: 0] regfile_out2;   // out2 of regfile

    wire    [ 4: 0] mux1_out;       // IF ID
    wire    [31: 0] mux2_out;       // ID EX
    wire    [31: 0] mux3_out;       // MEM WB
    wire    [31: 0] mux4_out;
    wire    [ 4: 0] mux5_out;
    wire    [31: 0] mux6_out;

    wire    [ 3: 0] alu_ctrl_out;   // out of alu controller
    wire    [31: 0] alu_out;        // out of alu
    wire    [31: 0] dm_out;         // out of dm
    wire    [31: 0] branch_add_out; // out of branch add

    // pipeline register
    wire  [31: 0] IF_ID_pc_add_out;
    wire  [31: 0] IF_ID_im_out;

    wire  [ 1: 0] ID_EX_LS_bit;  
    wire          ID_EX_RegDst;  
    wire  [ 1: 0] ID_EX_Branch;  
    wire          ID_EX_MemtoReg;
    wire  [ 3: 0] ID_EX_ALUOp;
    wire          ID_EX_MemWrite;
    wire          ID_EX_ALUSrc;
    wire          ID_EX_RegWrite;
    wire          ID_EX_Jump;
    wire          ID_EX_Ext_op;
    wire          ID_EX_PctoReg;
    wire  [31: 0] ID_EX_regfile_out1;
    wire  [31: 0] ID_EX_regfile_out2;
    wire  [31: 0] ID_EX_pc_add_out;
    wire  [25: 0] ID_EX_instr26;    

    wire  [ 1: 0] EX_MEM_LS_bit;        
    wire  [ 1: 0] EX_MEM_Branch;        
    wire          EX_MEM_MemtoReg;      
    wire          EX_MEM_MemWrite;      
    wire          EX_MEM_RegWrite;      
    wire          EX_MEM_Jump;
    wire          EX_MEM_Ext_op;        
    wire          EX_MEM_PctoReg;       
    wire  [31: 0] EX_MEM_branch_add_out;
    wire          EX_MEM_zero;
    wire  [31: 0] EX_MEM_pc_add_out;
    wire  [25: 0] EX_MEM_instr26;
    wire  [31: 0] EX_MEM_alu_out;
    wire  [31: 0] EX_MEM_regfile_out2;
    wire  [ 4: 0] EX_MEM_mux1_out;

    wire          MEM_WB_RegWrite;
    wire          MEM_WB_MemtoReg;
    wire          MEM_WB_PctoReg;
    wire  [31: 0] MEM_WB_pc_add_out;
    wire  [31: 0] MEM_WB_dm_out;
    wire  [31: 0] MEM_WB_alu_out;
    wire  [ 4: 0] MEM_WB_mux1_out;

    // pc module
    pc u_pc(
        .NPC(NPC),
        .clock(clock),
        .reset(reset),
        .PC(PC)
    );

    pc_add u_pc_add(
        .PC(PC),
        .pc_add_out(pc_add_out)
    );

    npc u_npc(
        .Jump(EX_MEM_Jump),
        .branch(EX_MEM_Branch),
        .zero(EX_MEM_zero),
        .EX_MEM_branch_add_out(EX_MEM_branch_add_out),
        .EX_MEM_pc_add_out(pc_add_out),
        .EX_MEM_instr26(EX_MEM_instr26),
        .NPC(NPC)
    );

    // IF module, from pc value to the cycle's instructions
    im_4k u_im_4k(
        .pc(PC),
        .out_instr(instruction)
    );

    // IF/ID 
    IF_ID u_IF_ID(
        .clock(clock),
        .pc_add_out(pc_add_out),
        .im_out(instruction),
        .IF_ID_pc_add_out(IF_ID_pc_add_out),
        .IF_ID_im_out(IF_ID_im_out)
    );

    // ID module
    regfile u_regfile(
        .rs(IF_ID_im_out[25:21]),
        .rt(IF_ID_im_out[20:16]),
        .rd(mux5_out),
        .data(mux4_out),
        .RegWrite(MEM_WB_RegWrite),
        .clock(clock),
        .reset(reset),
        .regfile_out1(regfile_out1),
        .regfile_out2(regfile_out2)
    );

    // ID/EX
    ID_EX u_ID_EX(
        .clock(clock),
        .reset(reset),

        .LS_bit(LS_bit),
        .RegDst(RegDst),
        .Branch(Branch),
        .MemtoReg(MemtoReg),
        .ALUOp(ALUOp),
        .MemWrite(MemWrite),
        .ALUSrc(ALUSrc),
        .RegWrite(RegWrite),
        .Jump(Jump),
        .Ext_op(Ext_op),
        .PctoReg(PctoReg),
        .IF_ID_pc_add_out(IF_ID_pc_add_out),
        .regfile_out1(regfile_out1),
        .regfile_out2(regfile_out2),
        .instr26(IF_ID_im_out[25:0]),

        .ID_EX_LS_bit(ID_EX_LS_bit),
        .ID_EX_RegDst(ID_EX_RegDst),   
        .ID_EX_Branch(ID_EX_Branch),
        .ID_EX_MemtoReg(ID_EX_MemtoReg),
        .ID_EX_ALUOp(ID_EX_ALUOp),
        .ID_EX_MemWrite(ID_EX_MemWrite),
        .ID_EX_ALUSrc(ID_EX_ALUSrc),
        .ID_EX_RegWrite(ID_EX_RegWrite),
        .ID_EX_Jump(ID_EX_Jump),
        .ID_EX_Ext_op(ID_EX_Ext_op),
        .ID_EX_PctoReg(ID_EX_PctoReg),
        .ID_EX_regfile_out1(ID_EX_regfile_out1),    
        .ID_EX_regfile_out2(ID_EX_regfile_out2),
        .ID_EX_pc_add_out(ID_EX_pc_add_out),
        .ID_EX_instr26(ID_EX_instr26)
    );

    // EX module
    mux1 u_mux1(
        .rt(ID_EX_instr26[20:16]),
        .rd(ID_EX_instr26[15:11]),
        .RegDst(ID_EX_RegDst),
        .DstReg(mux1_out)
    );

    Ext u_Ext(
        .input_num(ID_EX_instr26[15:0]),
        .Ext_op(ID_EX_Ext_op),
        .output_num(ext_out) 
    );

    alu_ctrl u_alu_ctrl(
        .funct(ext_out[5:0]),           // last 5 bit of instruction, which repersents funct code
        .ALUOp(ID_EX_ALUOp),            // ALUOp
        .alu_ctrl_out(alu_ctrl_out)
    );

    mux2 u_mux2(
        .out2(ID_EX_regfile_out2),        // regfile_out2
        .Ext(ext_out),
        .ALUSrc(ID_EX_ALUSrc),            // ALUSrc
        .DstData(mux2_out)
    );

    alu u_alu(
        .op_num1(ID_EX_regfile_out1),     // regfile_out1
        .op_num2(mux2_out),
        .shamt(ext_out[10:6]),  
        .alu_ctrl_out(alu_ctrl_out),
        .zero(zero),
        .alu_out(alu_out)
    );

    branch_add u_branch_add(
        .ID_EX_pc_add_out(ID_EX_pc_add_out),
        .Ext_out(ext_out),
        .branch_add_out(branch_add_out)
    );

    mux6 u_mux6(
        .ID_EX_pc_add_out(ID_EX_pc_add_out),
        .ID_EX_regfile_out1(ID_EX_regfile_out1),
        .funct(ID_EX_instr26[5:0]),
        .mux6_out(mux6_out)
    );  

    // EX/MEM
    EX_MEM u_EX_MEM(
        .clock(clock),
        .reset(reset),

        .LS_bit(LS_bit),
        .Branch(ID_EX_Branch),
        .MemtoReg(ID_EX_MemtoReg),
        .MemWrite(ID_EX_MemWrite),
        .RegWrite(ID_EX_RegWrite),
        .Jump(ID_EX_Jump),
        .Ext_op(ID_EX_Ext_op),
        .PctoReg(ID_EX_PctoReg),

        .branch_add_out(branch_add_out),
        .zero(zero),
        .ID_EX_pc_add_out(mux6_out),
        .ID_EX_instr26(ID_EX_instr26),
        .alu_out(alu_out),
        .ID_EX_regfile_out2(ID_EX_regfile_out2),
        .mux1_out(mux1_out),

        .EX_MEM_LS_bit(EX_MEM_LS_bit),
        .EX_MEM_Branch(EX_MEM_Branch),
        .EX_MEM_MemtoReg(EX_MEM_MemtoReg),
        .EX_MEM_MemWrite(EX_MEM_MemWrite),
        .EX_MEM_RegWrite(EX_MEM_RegWrite),
        .EX_MEM_Jump(EX_MEM_Jump),
        .EX_MEM_Ext_op(EX_MEM_Ext_op),
        .EX_MEM_PctoReg(EX_MEM_PctoReg),
        .EX_MEM_branch_add_out(EX_MEM_branch_add_out),
        .EX_MEM_zero(EX_MEM_zero),
        .EX_MEM_pc_add_out(EX_MEM_pc_add_out),
        .EX_MEM_instr26(EX_MEM_instr26),
        .EX_MEM_alu_out(EX_MEM_alu_out),
        .EX_MEM_regfile_out2(EX_MEM_regfile_out2),
        .EX_MEM_mux1_out(EX_MEM_mux1_out)
    );

    
    // MEM module
    dm_4k u_dm_4k(
        .clock(clock),
        .EX_MEM_alu_out(EX_MEM_alu_out),
        .EX_MEM_regfile_out2(EX_MEM_regfile_out2),
        .LS_bit(EX_MEM_LS_bit),
        .MemWrite(EX_MEM_MemWrite),
        .Ext_op(EX_MEM_Ext_op),
        .dm_out(dm_out)
    );

    // MEM/WB
    MEM_WB u_MEM_WB(
        .clock(clock),
        .reset(reset),

        .RegWrite(EX_MEM_RegWrite),
        .MemtoReg(EX_MEM_MemtoReg),
        .PctoReg(EX_MEM_PctoReg),

        .EX_MEM_pc_add_out(EX_MEM_pc_add_out),
        .dm_out(dm_out),
        .EX_MEM_alu_out(EX_MEM_alu_out),
        .EX_MEM_mux1_out(EX_MEM_mux1_out),

        .MEM_WB_RegWrite(MEM_WB_RegWrite),
        .MEM_WB_MemtoReg(MEM_WB_MemtoReg),
        .MEM_WB_PctoReg(MEM_WB_PctoReg),
        .MEM_WB_pc_add_out(MEM_WB_pc_add_out),
        .MEM_WB_dm_out(MEM_WB_dm_out),
        .MEM_WB_alu_out(MEM_WB_alu_out),
        .MEM_WB_mux1_out(MEM_WB_mux1_out)
    );

    // WB module
    mux3 u_mux3(
        .dm_out(MEM_WB_dm_out),
        .alu_out(MEM_WB_alu_out),
        .MemtoReg(MEM_WB_MemtoReg),
        .mux3_out(mux3_out)
    );


    mux4 u_mux4(
        .mux3_out(mux3_out),
        .MEM_WB_pc_add_out(MEM_WB_pc_add_out),
        .PctoReg(MEM_WB_PctoReg),
        .mux4_out(mux4_out)
    );

    mux5 u_mux5(
        .MEM_WB_mux1_out(MEM_WB_mux1_out),
        .PctoReg(PctoReg),
        .mux5_out(mux5_out)
    );

endmodule
