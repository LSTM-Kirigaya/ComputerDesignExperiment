// `include "v1.v"
// `include "v2.v"
// `include "v3.v"

module main;
    v1 u_v1();
    v2 u_v2();
    v3 u_v3();
endmodule