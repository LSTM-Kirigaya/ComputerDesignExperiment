module Cause (
    
);

endmodule //Cause