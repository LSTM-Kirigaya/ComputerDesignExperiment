`include "./Controller/controller.v"
`timescale 10ns/10ns

module controller_tb();
    

endmodule //controller_tb