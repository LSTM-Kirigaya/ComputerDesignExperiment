module controller(opcode, RegDst, Branch, MemtoReg, ALUOp, 
    MemWrite, ALUSrc, RegWrite, Jump, Ext_op);

    input      [ 5: 0] opcode;         // 6-bit opcode, which is instr[31:26]         
    
    // outputs are all signals
    output reg         RegDst;   
    output reg         Branch;
    output reg         MemtoReg;
    output reg [ 3: 0] ALUOp;
    output reg         MemWrite;
    output reg         ALUSrc;
    output reg         RegWrite;
    output reg         Jump;
    output reg         Ext_op;

    // for easy use 
    `define SIGNAL {RegDst, Branch, MemtoReg, ALUSrc, ALUOp, MemWrite, RegWrite, Jump, Ext_op}
    parameter T = 1'b1;
    parameter F = 1'b0;

    /* opcode field */
    parameter opcode_is_RType  = 6'b000000;

    // conditional transfer
    parameter opcode_is_BEQ    = 6'b000100;
    parameter opcode_is_BNE    = 6'b000101;

    // I type R op
    parameter opcode_is_ADDI   = 6'b001000;
    parameter opcode_is_ADDIU  = 6'b001001;
    parameter opcode_is_LUI    = 6'b001111;
    parameter opcode_is_ORI    = 6'b001101;
    parameter opcode_is_XORI   = 6'b001110;
    parameter opcode_is_SLTI   = 6'b001010;
    parameter opcode_is_SLTIU  = 6'b001011;

    // load and save
    parameter opcode_is_LW     = 6'b100011;
    parameter opcode_is_LH     = 6'b100001;
    parameter opcode_is_LHU    = 6'b100101;
    parameter opcode_is_LB     = 6'b100000;
    parameter opcode_is_LBU    = 6'b100100;
    parameter opcode_is_SW     = 6'b101011;
    parameter opcode_is_SH     = 6'b101001;
    parameter opcode_is_SB     = 6'b101000;

    // J Type
    parameter opcode_is_J      = 6'b000010;
    parameter opcode_is_JAL    = 6'b000011;

    always @(*) 
    begin
        if (opcode == opcode_is_RType)    // R type operation, use funct
            `SIGNAL = {T, F, F, F, 4'b0010, F, T, F, F};
        else
            case(opcode) 
                // About ALUOp of I type and J type:
                // 0000: use add
                // 0001: use minus
                // 0011: load to upper 16-bit
                // 0100: use or
                // 0110: use xor
                // 1000: use slt
                opcode_is_BEQ   : `SIGNAL = {F, T, F, F, 4'b0001, F, F, F, F};
                opcode_is_BNE   : `SIGNAL = {F, T, F, F, 4'b0001, F, F, F, F};

                opcode_is_ADDI  : `SIGNAL = {F, F, F, T, 4'b0000, F, T, F, F};
                opcode_is_ADDIU : `SIGNAL = {F, F, F, T, 4'b0000, F, T, F, T};
                opcode_is_LUI   : `SIGNAL = {F, F, F, T, 4'b0011, F, T, F, F};
                opcode_is_ORI   : `SIGNAL = {F, F, F, T, 4'b0100, F, T, F, F};
                opcode_is_XORI  : `SIGNAL = {F, F, F, T, 4'b0110, F, T, F, F};
                opcode_is_SLTI  : `SIGNAL = {F, F, F, T, 4'b1000, F, T, F, F};
                opcode_is_SLTIU : `SIGNAL = {F, F, F, T, 4'b1000, F, T, F, T};
                
                opcode_is_LW    : `SIGNAL = {F, F, T, T, 4'b0000, F, T, F, F};
                opcode_is_LH    : `SIGNAL = {F, F, T, T, 4'b0000, F, T, F, F};
                opcode_is_LHU   : `SIGNAL = {F, F, T, T, 4'b0000, F, T, F, T};
                opcode_is_LB    : `SIGNAL = {F, F, T, T, 4'b0000, F, T, F, F};
                opcode_is_LBU   : `SIGNAL = {F, F, T, T, 4'b0000, F, T, F, T};
                opcode_is_SW    : `SIGNAL = {F, F, F, T, 4'b0000, T, F, F, F};
                opcode_is_SH    : `SIGNAL = {F, F, F, T, 4'b0000, T, F, F, F};
                opcode_is_SB    : `SIGNAL = {F, F, F, T, 4'b0000, T, F, F, F};
    
                opcode_is_J     : `SIGNAL = {F, F, F, F, 4'b0000, F, F, T, F};
                opcode_is_JAL   : `SIGNAL = {F, F, F, F, 4'b0000, F, T, T, F};

            endcase    
    end
endmodule